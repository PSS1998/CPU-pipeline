module Datapath(input reset, clk, input sel_stack , input [1:0] PCsrc, input push, pop, RegDt, input [1:0] ALUsrc, input [2:0] ALUop, input shift, MemRead, MemWrite, MemtoReg, RegWrite, input change_zero_carry, output zero, carry, output const_sign, output[4:0] inst, output WB_RegWrite, MEM_RegWrite, output [2:0] MEM_RegRd, WB_RegRd, EX_RegRs, EX_RegRt, input[1:0] ForwardA, input[1:0] ForwardB, output EX_MemRead, output [2:0] EX_RegRd, output [2:0] ID_RegRs, output [2:0] ID_RegRt, output [5:0] inst2, input ldPC, input ld_IF_ID, input ID_EX_flush, input sel_carry_forwarding, sel_zero_forwarding, carry_forwarding, zero_forwarding, output logic [2:0] inst3, output logic EX_change_C_Z, zero_out, carry_out);
  
  logic[11:0] PC_in;
  logic[11:0] PC_out;
  logic[11:0] PC_plus;
  logic[11:0] PC_jmp;
  logic[11:0] PC_jc;
  logic[11:0] PC_Mux_out;
  logic[11:0] stack_out;
  logic[18:0] instruction;
  logic[18:0] ID_inst;
  logic[11:0] ID_PC;
  logic[2:0] WB_WriteReg;
  logic[2:0] Reg_src2;
  logic[7:0] Reg_WriteData;
  logic[7:0] Read1;
  logic[7:0] Read2;
  logic[11:0] address_se;
  logic[16:0] control_signals;
  logic[16:0] ID_control;
  logic[7:0] EX_read1;
  logic[7:0] EX_read2;
  logic[7:0] shift_count;
  logic[7:0] const_EX;
  logic[16:0] EX_control_signal;
  logic[7:0] EX_const_EX;
  logic[7:0] EX_shift_count;
  logic[2:0] EX_inst10_8;
  logic[2:0] EX_inst7_5;
  logic[2:0] EX_inst13_11;
  logic[3:0] EX_control_signal2;
  logic[7:0] ALU1;
  logic[7:0] ALU2;
  logic[7:0] ALUsrc2;
  logic[7:0] MEM_ALUout;
  logic[7:0] ALUout;
  logic[2:0] Reg_Rt;
  logic[3:0] MEM_control_signal;
  logic[7:0] MEM_read2;
  logic[7:0] readMem;
  logic[1:0] WB_control_signal;
  logic[7:0] WB_Read_data;
  logic[7:0] WB_ALU_result;
  logic[2:0] WB_register_num;
  logic carry1;
  logic zero1;
  
  assign control_signals = {sel_stack , PCsrc, push, pop, RegDt, ALUsrc, ALUop, shift, MemRead, MemWrite, MemtoReg, RegWrite, change_zero_carry};
  //tedad bit control signala ghalate
  assign inst = ID_inst[18:14];
  assign inst2 = ID_inst[18:13];
  assign inst3 = ID_inst[18:16];
//  assign EX_Flush = ID_EX_flush;
  assign WB_WriteReg = WB_RegRd;
  assign EX_MemRead = EX_control_signal[4];
  assign EX_RegRd = EX_inst13_11;
  assign EX_RegRt = EX_inst10_8;
  assign ID_RegRs = ID_inst[7:5];
  assign ID_RegRt = ID_inst[10:8];
  assign EX_RegRs = EX_inst7_5;
  assign WB_RegWrite = WB_control_signal[0];
  assign MEM_RegWrite = MEM_control_signal[0];
  assign EX_change_C_Z = EX_control_signal[0];
 
  reg1 _reg1 (reset, clk, ID_EX_flush, EX_Flush);
  
  PC _PC (reset, clk, ldPC, PC_in, PC_out);
  adderPC _adderPC (PC_out, PC_plus);
  Mux12_3to1 Mux_src (PC_plus, PC_jc, ID_inst[11:0], PCsrc, PC_Mux_out);
  Mux12_2to1 Mux_src_stack (PC_Mux_out, stack_out, sel_stack, PC_in);
  InstMem _InstMem (clk, PC_out, instruction);
  IF_ID_reg _IF_ID_reg (clk, ld_IF_ID, IF_Flush, instruction, PC_plus, ID_inst, ID_PC);
  Mux3_2to1 Mux_Register (ID_inst[7:5], ID_inst[13:11], RegDt, Reg_src2);
  Register_file _Register_file (clk, ID_inst[10:8], Reg_src2, WB_WriteReg, Reg_WriteData, WB_control_signal[0], Read1, Read2);
  Stack _Stack (clk, pop, push, ID_PC, stack_out);
  sign_extend_8to12 _sign_extend_8to12 (ID_inst[7:0], address_se);
  adder2 _adder2 (ID_PC, address_se, PC_jc);
  Mux10_2to1 Mux_EX_flush (control_signals, ID_EX_flush, ID_control);
  sign_extend3to8 _sign_extend3to8 (ID_inst[3:0], shift_count);
  ID_EX_reg _ID_EX_reg (clk, ID_control, Read1, Read2, ID_inst[7:0], shift_count, ID_inst[10:8], ID_inst[7:5], ID_inst[13:11], EX_control_signal, EX_read1, EX_read2, EX_const_EX, EX_shift_count, EX_inst10_8, EX_inst7_5, EX_inst13_11);
  Mux4_2to1 Mux_MEM_WB_flush (EX_control_signal[4:1], EX_Flush, EX_control_signal2);
  Mux8_3to1 _ForwardA (EX_read1, Reg_WriteData, MEM_ALUout, ForwardA, ALU1);
  Mux8_3to1 _ForwardB (EX_read2, Reg_WriteData, MEM_ALUout, ForwardB, ALU2);
  Mux8_3to1 Mux_ALUsrc2 (ALU2, EX_const_EX, EX_shift_count, EX_control_signal[10:9], ALUsrc2);
  ALU _ALU (clk, ALU1, ALUsrc2, carry, EX_control_signal[5], EX_control_signal[8:6], ALUout, zero_out, carry_out);
  C_FF _C_FF (reset, clk, carry_out, EX_control_signal[0] , carry1);
  Mux1_2to1 Mux_carry_forwarding (carry1, carry_forwarding, sel_carry_forwarding, carry);
  Z_FF _Z_FF (reset, clk, zero_out, EX_control_signal[0], zero1);
  Mux1_2to1 Mux_zero_forwarding (zero1, zero_forwarding, sel_zero_forwarding, zero);
  Mux3_2to1 Mux_RegRt(EX_inst10_8, EX_inst13_11, EX_control_signal[11], Reg_Rt);
  EX_MEM_reg _EX_MEM_reg (clk, EX_control_signal2, ALUout, ALU2, EX_inst13_11, MEM_control_signal, MEM_ALUout, MEM_read2, MEM_RegRd);
  DataMemory _DataMemory (clk, MEM_ALUout, MEM_read2, MEM_control_signal[3], MEM_control_signal[2], readMem);
  MEM_WB_reg _MEM_WB_reg (clk, MEM_control_signal[1:0], readMem, MEM_ALUout, MEM_RegRd, WB_control_signal, WB_Read_data, WB_ALU_result, WB_RegRd);
  Mux8_2to1 Mux_WB (WB_Read_data, WB_ALU_result, WB_control_signal[1], Reg_WriteData);
  
endmodule
