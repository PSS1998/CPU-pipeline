module adder2(input[11:0] A, B, output[11:0] S);
   
  assign S = A+B;
  
endmodule
