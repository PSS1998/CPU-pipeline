`timescale 1ns/1ns
module InstMem(input clk, input[11:0] PC, output[18:0] instruction);
  
  logic[18:0] rom [4095:0];
  
// test 2
/*      initial  
      begin  
                rom[0] = 19'b0000011100000000000;  
                rom[1] = 19'b0000000100000000000;  
                rom[2] = 19'b0101001100100010100;  
                rom[3] = 19'b1010000000000000110;  
                rom[4] = 19'b1000001000101100100;  
                rom[5] = 19'b0001001111101000000; 
                rom[6] = 19'b1011100000000000001;  
                rom[7] = 19'b0000011101000000000;  
                rom[8] = 19'b0100000100100000001;  
                rom[9] = 19'b1110000000000000010;  
                rom[10] = 19'b0000000000000000000;  
                rom[11] = 19'b0000000000000000000;  
                rom[12] = 19'b0000000000000000000;  
                rom[13] = 19'b0000000000000000000;  
                rom[14] = 19'b0000000000000000000;  
                rom[15] = 19'b0000000000000000000;  
      end  
*/
	  initial  
      begin  
                rom[0] = 19'b1000000100001100100;  
                rom[1] = 19'b1000001000001100110;  
                rom[2] = 19'b0000001100101000000;  
                rom[3] = 19'b1000101100001101000;  
                rom[4] = 19'b1000000100001100101;  
                rom[5] = 19'b1000001000001100111; 
                rom[6] = 19'b0000101100101000000;    
                rom[7] = 19'b1000101100001101001;  
      end 
	
      assign instruction = (PC[11:0] < 4096 )? rom[PC]: 19'b0;  
  

  
endmodule



