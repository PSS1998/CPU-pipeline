module adderPC(input[11:0] A, output[11:0] S);
   
  assign S = A+1;
  
endmodule







